LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY sync_count_16bit IS 
	GENERIC (N : integer:=16);
	PORT (SW : IN STD_LOGIC_VECTOR(1 DOWNTO 0);
			KEY : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
			HEX0 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX1 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX2 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0);
			HEX3 : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
			);
END sync_count_16bit;
			
ARCHITECTURE Structural OF sync_count_16bit IS
	COMPONENT sync_count_16bit_block
		PORT (INPUT  : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
				OUTPUT : OUT STD_LOGIC
			);
END COMPONENT;
	COMPONENT decoder
		PORT ( I_D : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
			 HEX : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
			);	
END COMPONENT;
SIGNAL  CLK, ENBL, CLR : STD_LOGIC;
SIGNAL Q : STD_LOGIC_VECTOR(N-1 DOWNTO 0);
BEGIN 
--ASSEGNAZIONI 
ENBL<=SW(1);
CLR<=SW(0);
CLK<=KEY(0);

	FF_0 : sync_count_16bit_block PORT MAP (INPUT(0)=>ENBL, INPUT(1)=>CLK, INPUT(2)=>CLR, OUTPUT=>Q(0));
Count_cycle : FOR i IN 1 TO N-1 GENERATE 
	FF : sync_count_16bit_block PORT MAP (INPUT(0)=>Q(i-1), INPUT(1)=>CLK, INPUT(2)=>CLR, OUTPUT=>Q(i));
	END GENERATE;
--DECODER 
HEX_0 : decoder PORT MAP (I_D=>Q(3 DOWNTO 0), HEX=>HEX0);
HEX_1 : decoder PORT MAP (I_D=>Q(7 DOWNTO 4), HEX=>HEX1);
HEX_2 : decoder PORT MAP (I_D=>Q(11 DOWNTO 8), HEX=>HEX2);
HEX_3 : decoder PORT MAP (I_D=>Q(15 DOWNTO 12), HEX=>HEX3);
END Structural;


